module test;

logic a;

endmodule
