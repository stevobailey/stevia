//////////////////////////////////////////////////////////////////////////////
//
// author: Stevo Bailey (stevo.bailey@gmail.com)
//
// AES package
//
//////////////////////////////////////////////////////////////////////////////

package stv_aes_pkg;

  typedef enum logic [1:0] {
    AES128,
    AES192,
    AES256
  } stv_aes_keylen_t;

endpackage : stv_aes_pkg

