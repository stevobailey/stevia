module test;

logic a;
logic b;

endmodule
